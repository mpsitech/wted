-- file Crc8005_8.vhd
-- Crc8005_8 crcspec_v3_0 implementation
-- copyright: (C) 2016-2020 MPSI Technologies GmbH
-- author: Alexander Wirthmueller (auto-generation)
-- date created: 30 Jun 2024
-- IP header --- ABOVE

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Crc8005_8 is
	generic (
		initOneNotZero: boolean := false
	);
	port (
		reset: in std_logic;
		mclk: in std_logic;

		AXIS_tready: out std_logic;
		AXIS_tvalid: in std_logic;
		AXIS_tdata: in std_logic_vector(7 downto 0);
		AXIS_tlast: in std_logic;

		crc: out std_logic_vector(15 downto 0);
		validCrc: out std_logic
	);
end Crc8005_8;

architecture Rtl of Crc8005_8 is

	------------------------------------------------------------------------
	-- signal declarations
	------------------------------------------------------------------------

	---- main operation (op)
	type stateOp_t is (
		stateOpInit,
		stateOpCapt
	);
	signal stateOp: stateOp_t := stateOpInit;

	signal crc_sig: std_logic_vector(15 downto 0);
	signal validCrc_sig: std_logic;

begin

	------------------------------------------------------------------------
	-- implementation: main operation (op)
	------------------------------------------------------------------------

	AXIS_tready <= '1' when stateOp=stateOpCapt else '0';

	crc <= crc_sig;
	validCrc <= validCrc_sig;
	
	process (reset, mclk, stateOp)
		variable first: boolean;

	begin
		if reset='1' then
			stateOp <= stateOpInit;

			if not initOneNotZero then
				crc_sig <= (others => '0');
			else
				crc_sig <= (others => '1');
			end if;
			validCrc_sig <= '0';

			first := true;

		elsif rising_edge(mclk) then
			if stateOp=stateOpInit then
				if AXIS_tlast='0' then
					if not initOneNotZero then
						crc_sig <= (others => '0');
					else
						crc_sig <= (others => '1');
					end if;
					validCrc_sig <= '0';

					first := true;

					stateOp <= stateOpCapt;
				end if;

			elsif stateOp=stateOpCapt then
				if AXIS_tvalid='1' and (first or validCrc_sig='1') then
					crc_sig(15) <= AXIS_tdata(7) xor AXIS_tdata(6) xor AXIS_tdata(5) xor AXIS_tdata(4) xor AXIS_tdata(3) xor AXIS_tdata(2) xor AXIS_tdata(1) xor AXIS_tdata(0) xor crc_sig(7) xor crc_sig(8) xor crc_sig(9) xor crc_sig(10) xor crc_sig(11) xor crc_sig(12) xor crc_sig(13) xor crc_sig(14) xor crc_sig(15);
					crc_sig(14) <= crc_sig(6);
					crc_sig(13) <= crc_sig(5);
					crc_sig(12) <= crc_sig(4);
					crc_sig(11) <= crc_sig(3);
					crc_sig(10) <= crc_sig(2);
					crc_sig(9) <= AXIS_tdata(7) xor crc_sig(1) xor crc_sig(15);
					crc_sig(8) <= AXIS_tdata(7) xor AXIS_tdata(6) xor crc_sig(0) xor crc_sig(14) xor crc_sig(15);
					crc_sig(7) <= AXIS_tdata(6) xor AXIS_tdata(5) xor crc_sig(13) xor crc_sig(14);
					crc_sig(6) <= AXIS_tdata(5) xor AXIS_tdata(4) xor crc_sig(12) xor crc_sig(13);
					crc_sig(5) <= AXIS_tdata(4) xor AXIS_tdata(3) xor crc_sig(11) xor crc_sig(12);
					crc_sig(4) <= AXIS_tdata(3) xor AXIS_tdata(2) xor crc_sig(10) xor crc_sig(11);
					crc_sig(3) <= AXIS_tdata(2) xor AXIS_tdata(1) xor crc_sig(9) xor crc_sig(10);
					crc_sig(2) <= AXIS_tdata(1) xor AXIS_tdata(0) xor crc_sig(8) xor crc_sig(9);
					crc_sig(1) <= AXIS_tdata(7) xor AXIS_tdata(6) xor AXIS_tdata(5) xor AXIS_tdata(4) xor AXIS_tdata(3) xor AXIS_tdata(2) xor AXIS_tdata(1) xor crc_sig(9) xor crc_sig(10) xor crc_sig(11) xor crc_sig(12) xor crc_sig(13) xor crc_sig(14) xor crc_sig(15);
					crc_sig(0) <= AXIS_tdata(7) xor AXIS_tdata(6) xor AXIS_tdata(5) xor AXIS_tdata(4) xor AXIS_tdata(3) xor AXIS_tdata(2) xor AXIS_tdata(1) xor AXIS_tdata(0) xor crc_sig(8) xor crc_sig(9) xor crc_sig(10) xor crc_sig(11) xor crc_sig(12) xor crc_sig(13) xor crc_sig(14) xor crc_sig(15);
					validCrc_sig <= '1';

					first := false;

					if AXIS_tlast='1' then
						stateOp <= stateOpInit;
					end if;
				end if;
			end if;
		end if;
	end process;

end Rtl;
